----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 12/06/2022 06:09:18 PM
-- Design Name: 
-- Module Name: mux_1 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity mux_1 is
    Port( a, b, sel: in STD_LOGIC;
          res: out STD_LOGIC);
end mux_1;

architecture Behavioral of mux_1 is

begin
    
    process(sel, a, b)
    begin
    
    if sel = '1' then
        res <= b;
    else
        res <= a;
    end if;
    end process;
        

end Behavioral;
